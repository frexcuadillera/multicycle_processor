library verilog;
use verilog.vl_types.all;
entity signext_tb is
end signext_tb;
