library verilog;
use verilog.vl_types.all;
entity controllert is
end controllert;
