library verilog;
use verilog.vl_types.all;
entity s12_tb is
end s12_tb;
