library verilog;
use verilog.vl_types.all;
entity mem_tb is
end mem_tb;
